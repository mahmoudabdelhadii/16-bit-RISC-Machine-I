`define MREAD 2'b01
`define MWRITE 2'b10

`define RESET 5'b00000
`define WImm 5'b00001
`define LA 5'b00101
`define LB 5'b00100
`define ALU 5'b00110
`define regW 5'b00111
`define IF1 5'b01000
`define readM2 5'b01001
`define writeMD 5'b01010
`define Mwrite 5'b01011
`define readM 5'b01100
`define SetADR 5'b01101
`define LBR 5'b01110
`define ALU2 5'b01111
`define IF2 5'b10000
`define updatePC 5'b11000
`define decode 5'b11100
`define HALT 5'b11111

module cpu(clk,reset, mem_addr, mem_cmd, read_data, write_data);
input clk, reset;
input [15:0] read_data;
output [15:0] write_data;
output [8:0] mem_addr;
output [1:0] mem_cmd;

wire [2:0] readAndwrite,opcode;
wire [1:0] shift, op;
wire [15:0] sximm8;
wire [15:0] sximm5;
wire [11:0] FSM_out;
wire [15:0] Ireg_out;
wire [8:0] dataAddress;

wire[2:0] Z_out;
wire N,V,Z;

wire load_pc, load_addr, load_ir, reset_pc, addr_sel;

wire [8:0] next_pc,PC, intoOne,afterDataAddress;

assign intoOne = PC + 1;

vDFFE #(16) Instruction_Register(.clk(clk), .en(load_ir), .in(read_data), .out(Ireg_out)) ;

Instruction_Dec ID1(.in(Ireg_out), .nsel(FSM_out[11:9]),	//inputs
					.opcode(opcode), .op(op),				//to state machine
					.shift(shift), .sximm8(sximm8), .sximm5(sximm5), .readOrWrite(readAndwrite));	//to Datapath

FSM stateMachine(.opcode(opcode),.op(op),.reset(reset),.out(FSM_out),.clk(clk),.mem_cmd(mem_cmd), .addr_sel(addr_sel),.load_pc(load_pc),.reset_pc(reset_pc),.load_addr(load_addr), .load_ir(load_ir),.Z_out(Z_out),.N(N),.V(V),.Z(Z));


datapath DP(.mdata(read_data), .sximm8(sximm8), .sximm5(sximm5), .PC(8'b0), .writenum(readAndwrite), .write(FSM_out[0]), 
			.readnum(readAndwrite), .clk(clk), .asel(FSM_out[3]), .bsel(FSM_out[4]), .vsel(FSM_out[4:3]), .loadb(FSM_out[6]), .loada(FSM_out[5]), .loadc(FSM_out[7]), .loads(FSM_out[8]), .shift(shift), .ALUop(FSM_out[6:5]), 
			.datapath_out(write_data), .Z_out(Z_out), .N(N), .V(V), .Z(Z));
			

MUX #(9) PCMUX(.a(9'b0),.b(intoOne), .sel(reset_pc),.out(next_pc));
//module MUX(a,b,sel,out)

vDFFE #(9) ProgramCounter(.clk(clk), .en(load_pc), .in(next_pc), .out(PC));
vDFFE #(9) DataAddress(.clk(clk), .en(load_addr), .in(write_data[8:0]), .out(dataAddress));
//module vDFFE(clk, en, in, out)

MUX #(9) memSelect(.a(PC), .b(dataAddress),.sel(addr_sel),.out(mem_addr));




endmodule
module Instruction_Dec(in, nsel, opcode, op, shift, sximm8, sximm5, readOrWrite);
input [15:0] in;
input [2:0] nsel;

output [1:0] op,shift;
reg [1:0] shift;
output [2:0] opcode;
output [15:0] sximm8; //specify datapath size
output [15:0] sximm5;
output [2:0] readOrWrite; //check wire/reg here - writenum and readnum

wire [2:0] rORw;


assign opcode = in[15:13];
assign op = in [12:11];
//assign shift = in[4:3];
assign sximm8 = {{8{in[7]}}, in [7:0] };
assign sximm5 = {{11{in[4]}}, in [4:0] };
assign readOrWrite = rORw;

always @(*)
if (opcode == 3'b110 || opcode == 3'b101)
	shift = in[4:3];
else
	shift = 2'b00;


writeAndRead_Mux M1(.Rn(in[10:8]),.Rd(in[7:5]),.Rm(in[2:0]), .nsel(nsel),.readOrWrite(rORw) );


endmodule

module writeAndRead_Mux(Rn, Rd, Rm, nsel, readOrWrite);
input [2:0] Rn, Rd, Rm, nsel;

output [2:0] readOrWrite;

reg [2:0] readOrWrite;

always@*begin
	case(nsel)
		3'b001: readOrWrite = Rn;
		3'b010: readOrWrite = Rd;
		3'b100: readOrWrite = Rm;
		default: readOrWrite = 3'bxxx;
		
		//continue those
	endcase
end
endmodule





module FSM(opcode,op,reset,out,clk,mem_cmd, addr_sel,load_pc,reset_pc, load_addr, load_ir,Z_out,N,V,Z);
input clk;
input[2:0] opcode;
input[1:0] op;
input reset;

input [2:0] Z_out;
input N,V,Z;

output[11:0] out;
output addr_sel,load_pc,reset_pc,load_addr, load_ir;
output [1:0] mem_cmd;

reg[11:0] out;
reg addr_sel,load_pc,reset_pc,load_addr, load_ir;
reg [1:0] mem_cmd;

reg[4:0] state;

always@ (posedge clk) begin
	
	casex ({state,reset,opcode,op})
		
		//reset
		11'bxxxxx_1_xxx_xx : state = `reset; //reset state is still 00000
		
		//reset stage
		{`reset,6'b0_xxx_xx} : state = `IF1;	//advance to IF1

		//state 01000 IF1
		{`IF1,6'b0_xxx_xx} : state = `IF2;	//advance to IF2

		//state 10000 IF2
		{`IF2,6'b0_xxx_xx} : state = `updatePC;	//advance to UpdatePC

		//state 11000 UpdatePC
		{`updatePC,6'b0_xxx_xx} : state = `decode;	//advance to decode
		
		//state 11100 decode
		{`decode,6'b0_110_10} : state = `WImm;	//MOV Rn,#<im8>
		{`decode,6'b0_110_00} : state = `LB;	//MOV Rd,Rm{,<sh_op>}
		{`decode,6'b0_101_xx} : state = `LB;	//ALU instructions
		{`decode,6'b0_011_00} : state = `LA;	//LDR
		{`decode,6'b0_100_00} : state = `LA;	//STR
		{`decode,6'b0_111_xx} : state = `HALT;	//HALT
		//  ^^^ changed them to start taking messages from the decode state

		//state 00100 Load B
		{`LB,6'b0_101_0x} : state = `LA;	//Load A
		{`LB,6'b0_101_10} : state = `LA;	//Load A 
		{`LB,6'b0_110_00} : state = `ALU;	//ALU
		{`LB,6'b0_101_11} : state = `ALU;	//ALU

		//state 00001 writeImm
		{`WImm,6'b0_xxx_xx} : state = `IF1; 	//IF1
		
		//state 00101 Load A
		{`LA,6'b0_xxx_xx : state} = `ALU;	//always goes to ALU
		
		//state 00110 ALU operations
		{`ALU,6'b0_101_01} : state = `IF1;	//CMP - IF1
		{`ALU,6'b0_110_00} : state =`IF1;	//IF1
		{`ALU,6'b0_101_00} : state = `IF1;	//IF1
		{`ALU,6'b0_101_1x} : state = `IF1;	//IF1
		{`ALU,6'b0_011_00} : state = `readM;	//LDR - ReadMem
		{`ALU,6'b0_100_00} : state = `setADR;	//STR - SetARD
		
		//state 00111 writeReg
		{`regW,6'b0_xxx_xx} : state = `IF1;
		
		//state 01100 readMem (LDR)
		{`readM,6'b0_xxx_xx} : state = `readM2;	//always goes to writeMD
		
		//state 01001 readMem2 (LDR)
		{`readM2,6'b0_xxx_xx} : state = `writeMD;
		
		//state 01010 WriteMD (LDR)
		{`writeMD,6'b00_xxx_xx} : state = `IF1;	//always goes to IF1
		
		//state 01101 SetADR (STR)
		{`setADR,6'b0_xxx_xx} : state = `LBR;	//always goes to LoadBR
		
		//state 01110 LoadBR (STR)
		{`LBR,6'b0_xxx_xx} : state = `ALU2;	//always goes to ALU2
		
		//state 01111 ALU2 (STR)
		{`ALU2,6'b0_xxx_xx} : state = `Mwrite;	//always goes to Mwrite
		
		//state 01011 Mwrite (STR)
		{`Mwrite,6'b0_xxx_xx} : state = `IF1;	//always goes to IF1

		//state 11111 HALT
		{`HALT,6'b0_xxx_xx} : state = `HALT;
		
		default : state = 5'bxxxxx;
	endcase
	
	case (state)

		//reset
		`reset : begin 
		out = 12'b000_00000000_0;
			//w = 2'b01;
		reset_pc = 1;
		load_pc  = 1;
		end
		
		//IF1
		`IF1 : begin
		out = 12'b000_00000000_0;
		reset_pc = 0;
		load_pc = 0;
		addr_sel = 1;
		mem_cmd = `MREAD;
		end
		
		//IF2
		`IF2 : begin
		addr_sel = 1;
		mem_cmd = `MREAD;
		load_ir = 1;
		end

		//Update PC
		`updatePC : begin
		mem_cmd = 2'b0;
		load_ir = 0;
		load_pc = 1;
		end

		//Decode
		`decode : begin
			load_pc = 0;
			out = 12'b0000000_11_000;	//defaults selects to 1
		end
		
		//writeImm
		`WImm : begin
			out = 12'b001_0000_10_00_1;
		end
		
		//loadB
		`LB : begin
			out = {(7'b100_0010), 2'b01, (3'b0)};
		end
		
		//loadA
		`LA : out = {(7'b001_0001),out[4], 1'b0, (3'b0)};
		
		//ALU instructions
		`ALU : out = {3'b000_,({opcode,op}==5'b10101 ? 1 : 0),1'b1,op,out[4],out[3],3'b00_0};
	
		//writeReg
		`regW : out = 12'b010_00000000_1;
		
		//readMem
		5'b01100: begin
		`readM = 1; addr_sel = 0; mem_cmd = `MREAD;
		end
		
		//readMem2
		`readM2 : begin
		end
		
		//writeMD
		`writeMD : begin
		out = 12'b010_000011001;
		end
		
		//SetADR
		`setADR : begin
		load_addr = 1; addr_sel = 0;
		end
		
		//LoadBR
		`LBR : begin
		out = {(7'b010_0010), 2'b01, (3'b0)};
		end
		
		//ALU2
		`ALU2 : begin
		out = {5'b000_01,op,out[4],out[3],3'b00_0};
		end
		
		//Mwrite
		`Mwrite : begin
		mem_cmd = `MWRITE;
		end
		
		//HALT
		`HALT : begin
		end
		
		default : out = 12'b000000000000;
		
			
		
	endcase
	
	
end

endmodule







